module FPCVT(D, S, E, F);

   input wire [11:0] D;

   output reg        S;
   output reg [2:0]  E;
   output reg [3:0]  F;

   

endmodule
