module exp(D, E);

   input wire [10:0] mag;
   output wire [2:0] E;

   integer           i;
   
   always @(*) begin
      for (i = 0; i < 8; i = i + 1) begin
         
      end
   end

endmodule
