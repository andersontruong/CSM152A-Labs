module lze();


endmodule; // lze
