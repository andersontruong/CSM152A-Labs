module lze(a, q);

    input wire [1:0] a;
    output wire q;

    assign q = a[0];

endmodule; // lze
